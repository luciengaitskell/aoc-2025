// rtl/top.sv
module top (
    input clk,
    output logic out
);
  assign out = clk;
endmodule
